module mux2_1(s, d0, d1)



endmodule